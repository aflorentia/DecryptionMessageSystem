library verilog;
use verilog.vl_types.all;
entity samtest is
end samtest;
